`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 05/05/2023 12:19:19 PM
// Design Name: 
// Module Name: Mux3x1
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module Mux3x1(
 input read_data1IDEX,
 input [1:0] forward,
 input [4:0] result,
 input [4:0] rdEXMEM,
 input [4:0] rdMEMWB
    );
    
endmodule
